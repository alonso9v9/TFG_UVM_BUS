// Curso: EL-5617 Trabajo final de graduación
// Tecnologico de Costa Rica (www.tec.ac.cr)
// Desarrollador:
// Alonso Vega-Badilla (alonso_v_@estudiantec.cr)
// Este script esta estructurado en System Verilog
// Proposito General:
// Pacquete de parámetros


package bus_parameters;

    parameter pckg_sz=16;
    parameter drvrs=4;
    parameter fif_Size=10;
    parameter bits =16;

endpackage:bus_parameters